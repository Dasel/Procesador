----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:30:05 04/16/2016 
-- Design Name: 
-- Module Name:    adder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity adder is
		Port ( op1 : in  STD_LOGIC_VECTOR (31 downto 0);
				 op2 : in  STD_LOGIC_VECTOR (31 downto 0);
				 resultado : out  STD_LOGIC_VECTOR (31 downto 0));
end adder;

architecture arqAdder of adder is

begin
		process(op1,op2)
			begin
				resultado <= op1 + op2;
			end process;


end arqAdder;

